module UART_tx(input clk, input rst_n, output TX, input trmt, input [7:0] tx_data, output logic tx_done);

typedef enum logic {IDLE, CNT} state_t;
state_t state, nxt_state;
logic [8:0] tx_shft_reg;
logic init, shift, set_done,transmitting;
logic [11:0] baud_cnt;
logic [3:0] bit_cnt;

// TX data shifter
always_ff @(posedge clk, negedge rst_n)
	if (!rst_n)
		tx_shft_reg <= 9'h1ff;
	else if (init == 1'b1)
		tx_shft_reg <= {tx_data, 1'b0};
	else if (shift == 1'b1)
		tx_shft_reg <= {1'b1, tx_shft_reg[8:1]};

// baud counter 	
always_ff @(posedge clk, negedge rst_n)
	if (!rst_n)
		baud_cnt <= 12'h000;
	else if (init|shift == 1'b1)
		baud_cnt <= 12'h000;
	else if ({init|shift, transmitting} == 2'b01)
		baud_cnt <= baud_cnt +1;

// check if we have reach the hold period
assign shift = baud_cnt == 12'd2604;

// shift counter
always_ff @(posedge clk, negedge rst_n)
	if (!rst_n)
		bit_cnt <= 4'h0;
	else if (init == 1'b1)
		bit_cnt <= 4'h0;
	else if (shift == 1'b1)
		bit_cnt <= bit_cnt + 1;

// RS flop
always_ff @(posedge clk, negedge rst_n)
	if (!rst_n)
		tx_done <= 1'b0;
	else if (init)
		tx_done <= 1'b0;
	else if (set_done) 
		tx_done <= 1'b1;

// FSM flop
always_ff @(posedge clk, negedge rst_n)
	if (!rst_n)
		state <= IDLE;
	else 
		state <= nxt_state;

always_comb begin
	// initialize outputs to avoid latches
	init = 0;
	transmitting = 0;
	set_done = 0;
	nxt_state = state;

	case(state)
		default:
			if (trmt) begin
				init = 1'b1;
				state = CNT;
			end
		CNT:
			if (!bit_cnt != 4'd10) begin
				transmitting = 1'b1;
			end else begin
				set_done = 1'b1;
				nxt_state = IDLE;
			end
	endcase
end
endmodule