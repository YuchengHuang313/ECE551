module SDiv_tb();



endmodule
